module top (
    input  wire clk,            // system clock
    input  wire rst_n,          // active low reset
    input  wire rx,             // from STM32 TX

    output wire [6:0] seg_tens, // left 7-seg (high digit)
    output wire [6:0] seg_ones  // right 7-seg (low digit)
);

    // UART receiver
    wire [7:0] rx_byte;
    wire       rx_done;

    uart_rx #(
        .CLKS_PER_BIT(16)       // set according to your clock (10MHz -> 87)
    ) u_rx (
        .clk     (clk),
        .rst_n   (rst_n),
        .rx      (rx),
        .rx_byte (rx_byte),
        .rx_done (rx_done)
    );

    // BCD digits for two 7-seg displays
    reg [3:0] bcd_tens;
    reg [3:0] bcd_ones;

    
	
// �ݴ��һ�������ַ�
	reg       have_first;     // 0 = ��û�е�һλ��1 = �Ѿ��յ���һλ
	reg [7:0] first_ascii;    // �����һλ ASCII

	always @(posedge clk or negedge rst_n) begin
		 if (!rst_n) begin
			  bcd_tens   <= 4'd0;
			  bcd_ones   <= 4'd0;
			  have_first <= 1'b0;
			  first_ascii <= 8'd0;
		 end else begin
			  if (rx_done) begin
					// ֻ���� '0'..'9'�������ֽ�ֱ������
					if (rx_byte >= "0" && rx_byte <= "9") begin
						 if (!have_first) begin
							  // ������һ����ĵ�һλ����
							  first_ascii <= rx_byte;
							  have_first  <= 1'b1;
						 end else begin
							  // ���ǵڶ�λ���֣����һ�ԣ�first_ascii + rx_byte
							  bcd_tens   <= first_ascii - "0";  // ��λ
							  bcd_ones   <= rx_byte     - "0";  // ��λ
							  have_first <= 1'b0;               // ׼����һ��
						 end
					end
					// ������� '0'..'9' ����ȫ���ӣ����� bcd_tens / bcd_ones
			  end
		 end
	end
    bcd_to_seg u_seg_tens (
        .bcd (bcd_tens),
        .seg (seg_tens)
    );

    bcd_to_seg u_seg_ones (
        .bcd (bcd_ones),
        .seg (seg_ones)
    );

    // ������õ��ǹ�����������ܣ�������������һ��ȡ����
     wire [6:0] seg_tens_n = ~seg_tens;
     wire [6:0] seg_ones_n = ~seg_ones;
    // Ȼ���� UCF ��Լ�� seg_tens_n / seg_ones_n ��Ӧ���š�

endmodule
