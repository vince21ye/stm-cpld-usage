module shift_register_sipo #(
    parameter WIDTH = 8    // ��λ�Ĵ���λ���ɵ�
)(
    input  wire clk,       // ʱ��
    input  wire rst,       // ͬ����λ������Ч��
    input  wire shift_en,  // ��λʹ�ܣ�����Ч��
    input  wire serial_in, // �������� bit
    output reg  [WIDTH-1:0] parallel_out // ��������Ĵ���
);

    always @(posedge clk) begin
        if (rst) begin
            parallel_out <= {WIDTH{1'b0}};   // resest
        end 
        else if (shift_en) begin
            // The serial bit enters the most significant bit (MSB), and all other data shift right by one position.
            parallel_out <= {serial_in, parallel_out[WIDTH-1:1]};
        end
    end

endmodule
